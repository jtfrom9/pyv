module hoge;

endmodule

