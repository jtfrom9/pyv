module hoge()

endmodule

