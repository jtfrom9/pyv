module hoge(a,b,foo,bar)

endmodule

